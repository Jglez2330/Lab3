module notA_N #(parameter N = 8)
					(input logic[N-1:0] a, output logic[N-1:0] y);
					
					
		assign y = ~ a;
		

endmodule

