//Módulo AND de 3 bits


module and_3 (input logic H,J,K, output logic V);


			assign V = H & J & K;
			
			
endmodule