module AdderNBits #(parameter NBITS = 4)(input logic [NBITS-1 : 0] A, 
														input logic [NBITS-1 : 0] B,
														input logic Cin,
														output logic Cout,
														output logic [NBITS-1 : 0] result);


endmodule 