//Módulo XOR de 2 bits


module xor_2 (input logic yn1,an1, output logic J);


			assign J = yn1 ^ an1;
			
			
endmodule

