//Módulo XNOR de 2 bits


module xnor_2 (input logic an1,bn1, output logic K);


			assign J = ~(an1 ^ bn1);
			
			
endmodule
